module main;
  initial
    begin
      $display("Merry Christmas everybody !!");
      $finish ;
    end
endmodule